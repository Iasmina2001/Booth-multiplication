library verilog;
use verilog.vl_types.all;
entity booth_tb is
end booth_tb;
